library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;

entity ramtest is
	port(
		signal ram_type0 :  unsigned(15 downto 0) ;
		signal ram_type1 :  unsigned(15 downto 0) ;
		signal ram_type2 :  unsigned(15 downto 0) ;
		signal ram_type3 :  unsigned(15 downto 0) ;
		signal ram_type4 :  unsigned(15 downto 0) ;
		signal ram_type5 :  unsigned(15 downto 0) ;
		signal ram_type6 :  unsigned(15 downto 0) ;
		signal ram_type7 :  unsigned(15 downto 0) ;
		signal ram_type8 :  unsigned(15 downto 0) ;
		signal ram_type9 :  unsigned(15 downto 0) ;
		signal ram_type10 :  unsigned(15 downto 0) ;
		signal ram_type11 :  unsigned(15 downto 0) ;
		signal ram_type12 :  unsigned(15 downto 0) ;
		signal ram_type13 :  unsigned(15 downto 0) ;
		signal ram_type14 :  unsigned(15 downto 0) ;
		signal ram_type15 :  unsigned(15 downto 0) 
	);

end ramtest;

architecture rt of ramtest is
begin
end rt;
