-- Implements a simple Nios II system for the DE-series board.
-- Inputs: SW7-0 are parallel port inputs to the Nios II system
-- CLOCK_50 is the system clock
-- KEY0 is the active-low system reset
-- Outputs: LEDG7-0 are parallel port outputs from the Nios II system

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;

ENTITY integration IS
	PORT (
		SW : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		KEY : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		
		CLOCK_50 : IN STD_LOGIC;
		
		LEDG : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		DRAM_CLK, DRAM_CKE : OUT STD_LOGIC;
		DRAM_ADDR : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
		DRAM_BA_0, DRAM_BA_1 : BUFFER STD_LOGIC;
		DRAM_CS_N, DRAM_CAS_N, DRAM_RAS_N, DRAM_WE_N : OUT STD_LOGIC;
		DRAM_DQ : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		DRAM_UDQM, DRAM_LDQM : BUFFER STD_LOGIC;
		
		LCD_DATA : inout STD_LOGIC_VECTOR (7 downto 0);
		LCD_ON, LCD_BLON, LCD_EN, LCD_RW, LCD_RS : out STD_LOGIC;
		
		VGA_R:out	std_logic_vector(9	downto	0);	
		VGA_G:out	std_logic_vector(9	downto	0);	
		VGA_B:out	std_logic_vector(9	downto	0);	
		VGA_CLK:	out	std_logic;
		VGA_BLANK:	out	std_logic;	
		VGA_HS:out	std_logic;	
		VGA_VS:out	std_logic;	
		VGA_SYNC:out	std_logic;
		
		SRAM_DQ	:	INOUT	STD_LOGIC_VECTOR(15	downto	0);
		SRAM_ADDR	:	OUT	STD_LOGIC_VECTOR(17	downto	0);
		SRAM_LB_N	:	OUT	STD_LOGIC;
		SRAM_UB_N	:	OUT	STD_LOGIC;
		SRAM_CE_N	:	OUT	STD_LOGIC;
		SRAM_OE_N	:	OUT	STD_LOGIC;
		SRAM_WE_N	:	OUT	STD_LOGIC;
		
		SD_DAT, SD_DAT3, SD_CMD : inout std_LOGIC;
		SD_CLK : OUT STD_LOGIC;
		
		PS2_CLK		:	INOUT	STD_LOGIC;
		PS2_DAT		:	INOUT	STD_LOGIC;
		
		I2C_SDAT: inout STD_LOGIC;
		I2C_SCLK: OUT STD_LOGIC;
		AUD_XCK: OUT STD_LOGIC;
		CLOCK_27: IN STD_LOGIC;
		AUD_ADCDAT: IN STD_LOGIC;
		AUD_ADCLRCK: IN STD_LOGIC;
		AUD_BCLK: IN STD_LOGIC;
		AUD_DACDAT: inout STD_LOGIC;
		AUD_DACLRCK: IN STD_LOGIC);
END integration;

ARCHITECTURE Structure OF integration IS
COMPONENT nios_system
	PORT (
		clk_clk : IN STD_LOGIC;
		reset_reset_n : IN STD_LOGIC;
		sdram_clk_clk : OUT STD_LOGIC;
		
		key1_export : IN STD_LOGIC;
		key2_export : IN STD_LOGIC;
		key3_export : IN STD_LOGIC;
		
		leds_export : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		switches_export : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		
		sdram_wire_addr : OUT STD_LOGIC_VECTOR(11 DOWNTO 0);
		sdram_wire_ba : BUFFER STD_LOGIC_VECTOR(1 DOWNTO 0);
		sdram_wire_cas_n : OUT STD_LOGIC;
		sdram_wire_cke : OUT STD_LOGIC;
		sdram_wire_cs_n : OUT STD_LOGIC;
		sdram_wire_dq : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
		sdram_wire_dqm : BUFFER STD_LOGIC_VECTOR(1 DOWNTO 0);
		sdram_wire_ras_n : OUT STD_LOGIC;
		sdram_wire_we_n : OUT STD_LOGIC;

		-------------LCD--------------------
		lcd_data_DATA    : inout std_logic_vector(7 downto 0); --   lcd_data.DATA
		lcd_data_ON      : out   std_logic;                                        --           .ON
		lcd_data_BLON    : out   std_logic;                                        --           .BLON
		lcd_data_EN      : out   std_logic;                                        --           .EN
		lcd_data_RS      : out   std_logic;                                        --           .RS
		lcd_data_RW      : out   std_logic;                                        --           .RW

		-------------VGA--------------------
		vga_controller_CLK	: out std_logic;
		vga_controller_HS		: out std_logic;
		vga_controller_VS		: out std_logic;
		vga_controller_BLANK : out std_logic;
		vga_controller_SYNC	: out std_logic;
		vga_controller_R		: out std_logic_vector (9 downto 0);
		vga_controller_G		: out std_logic_vector (9 downto 0);
		vga_controller_B		: out std_logic_vector (9 downto 0);
		
		sram_DQ					: inout std_logic_vector (15 downto 0);
		sram_ADDR				: out std_logic_vector (17 downto 0);
		sram_LB_N				: out std_logic;
		sram_UB_N				: out std_logic;
		sram_CE_N				: out std_logic;
		sram_OE_N				: out std_logic;
		sram_WE_N				: out std_logic;
		
		-------------KEYBOARD---------------------
		ps2_keyboard_CLK		: inout std_logic;
		ps2_keyboard_DAT		: inout std_logic;

		clocks_clk_in_secondary_clk: IN STD_LOGIC;
		clocks_audio_clk_clk: out STD_LOGIC;
		
		sd_card_b_SD_dat : inout std_LOGIC;
		sd_card_b_SD_dat3 : inout std_LOGIC;
		sd_card_b_SD_cmd : inout std_LOGIC;
		sd_card_o_SD_clock : out std_LOGIC;
		
		audio_vid_SDAT: INOUT STD_LOGIC;
		audio_vid_SCLK: out STD_LOGIC;
		audio_ADCDAT: IN STD_LOGIC;
		audio_ADCLRCK: IN STD_LOGIC;
		audio_BCLK: IN STD_LOGIC;
		audio_DACDAT: out STD_LOGIC;
		audio_DACLRCK: IN STD_LOGIC);
END COMPONENT;

	SIGNAL DQM : STD_LOGIC_VECTOR(1 DOWNTO 0);
	SIGNAL BA : STD_LOGIC_VECTOR(1 DOWNTO 0);
	
BEGIN
	DRAM_BA_0 <= BA(0);
	DRAM_BA_1 <= BA(1);
	DRAM_UDQM <= DQM(1);
	DRAM_LDQM <= DQM(0);
--Instantiate the Nios II system entity generated by the Qsys tool.
	NiosII: nios_system
		PORT MAP (
			clk_clk => CLOCK_50,
			reset_reset_n => KEY(0),
			
			sdram_clk_clk => DRAM_CLK,
			
			leds_export => LEDG,
			
			key1_export => KEY(1),
			key2_export => KEY(2),
			key3_export => KEY(3),
			
			switches_export => SW,
			
			sdram_wire_addr => DRAM_ADDR,
			sdram_wire_ba => BA,
			sdram_wire_cas_n => DRAM_CAS_N,
			sdram_wire_cke => DRAM_CKE,
			sdram_wire_cs_n => DRAM_CS_N,
			sdram_wire_dq => DRAM_DQ,
			sdram_wire_dqm => DQM,
			sdram_wire_ras_n => DRAM_RAS_N,
			sdram_wire_we_n => DRAM_WE_N,
			
			lcd_data_DATA => LCD_DATA,
			lcd_data_ON => LCD_ON,
			lcd_data_BLON => LCD_BLON,
			lcd_data_EN => LCD_EN,
			lcd_data_RS => LCD_RS,
			lcd_data_RW => LCD_RW,
			
			vga_controller_CLK	=>	VGA_CLK,	
			vga_controller_HS	=>	VGA_HS,	
			vga_controller_VS	=>	VGA_VS,	
			vga_controller_BLANK	=>	VGA_BLANK,	
			vga_controller_SYNC	=>	VGA_SYNC,	
			vga_controller_R	=>	VGA_R,	
			vga_controller_G	=>	VGA_G,	
			vga_controller_B	=>	VGA_B,
			
			sram_DQ	=>	SRAM_DQ,
			sram_ADDR	=>	SRAM_ADDR,
			sram_LB_N	=>	SRAM_LB_N,
			sram_UB_N	=>	SRAM_UB_N,		
			sram_CE_N	=>	SRAM_CE_N,
			sram_OE_N	=>	SRAM_OE_N,
			sram_WE_N	=>	SRAM_WE_N,
		
			sd_card_b_SD_dat => SD_DAT,
			sd_card_b_SD_dat3 => SD_DAT3,
			sd_card_b_SD_cmd => SD_CMD,
			sd_card_o_SD_clock => SD_CLK,

			audio_vid_SDAT => I2C_SDAT,
			audio_vid_SCLK => I2C_SCLK,
			clocks_audio_clk_clk => AUD_XCK,
			clocks_clk_in_secondary_clk => CLOCK_27,
			audio_ADCDAT => AUD_ADCDAT,
			audio_ADCLRCK => AUD_ADCLRCK,
			audio_BCLK => AUD_BCLK,
			audio_DACDAT => AUD_DACDAT,
			audio_DACLRCK => AUD_DACLRCK,
			
			ps2_keyboard_CLK => PS2_CLK,
			ps2_keyboard_DAT => PS2_DAT);
	END Structure;